module ifu(
    input clk,
    input [31:0] pc,
    output [31:0] s
);
    

endmodule

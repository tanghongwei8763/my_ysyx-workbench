module ysyx_25020037_IFU(
    input clk,
    input [31:0] pc,
    output [31:0] s
);


endmodule
